�cclan
Clan
q.